library verilog;
use verilog.vl_types.all;
entity controlador_vertical1_vlg_vec_tst is
end controlador_vertical1_vlg_vec_tst;
